-- Name: DES_def.vhd
-- Author: Terry Huang
-- Description:
-- DES module permutaion, substitute table definition and some function
LIBRARY IEEE;
    USE IEEE.std_logic_1164.all;
    USE IEEE.std_logic_unsigned.all;
    USE IEEE.numeric_std.all;

PACKAGE DES_def IS
    -- Data definition
    SUBTYPE shift_Size IS integer range 0 to 2;
    SUBTYPE sel_Size IS integer range 0 to 15;
    SUBTYPE half_Size IS integer range 1 to 32;
    SUBTYPE key_Size IS integer range 1 to 56;
    SUBTYPE Size IS integer range 1 to 64;
    
    TYPE Init_Table IS ARRAY( 1 to 64 ) OF Size;
    TYPE PChoice_Table IS ARRAY( 1 to 28 ) OF Size;
    TYPE Expan_Table IS ARRAY( 1 to 48 ) OF half_Size;
    TYPE Permu_Table IS ARRAY( 1 to 32 ) OF half_Size;
    TYPE Permu_Sec_Table IS ARRAY( 1 to 48 ) OF key_Size;
    TYPE Box IS ARRAY( 0 to 3, 0 to 15) OF sel_Size;
    TYPE S_Box IS ARRAY( 1 to 8 ) OF Box;
    TYPE Shift_Table IS ARRAY( 1 to 17 ) OF shift_Size;

    Constant IP_Table : Init_Table := ( 58, 50, 42, 34, 26, 18, 10, 2,
                                        60, 52, 44, 36, 28, 20, 12, 4,
                                        62, 54, 46, 38, 30, 22, 14, 6,
                                        64, 56, 48, 40, 32, 24, 16, 8,
                                        57, 49, 41, 33, 25, 17,  9, 1,
                                        59, 51, 43, 35, 27, 19, 11, 3,
                                        61, 53, 45, 37, 29, 21, 13, 5,
                                        63, 55, 47, 39, 31, 23, 15, 7 );

    Constant IP_Inv_Table : Init_Table := ( 40, 8, 48, 16, 56, 24, 64, 32,
                                            39, 7, 47, 15, 55, 23, 63, 31,
                                            38, 6, 46, 14, 54, 22, 62, 30,
                                            37, 5, 45, 13, 53, 21, 61, 29,
                                            36, 4, 44, 12, 52, 20, 60, 28,
                                            35, 3, 43, 11, 51, 19, 59, 27,
                                            34, 2, 42, 10, 50, 18, 58, 26,
                                            33, 1, 41,  9, 49, 17, 57, 25 );
    
    Constant E_Table : Expan_Table := ( 32,  1,  2,	 3,	 4,	 5,
                                         4,  5,  6,	 7,	 8,	 9,
                                         8,  9, 10,	11,	12,	13,
                                        12, 13, 14,	15,	16,	17,
                                        16, 17,	18,	19,	20,	21,
                                        20, 21,	22,	23,	24,	25,
                                        24, 25,	26,	27,	28,	29,
                                        28, 29,	30,	31,	32,	 1 );

    Constant P_Table : Permu_Table := ( 16,  7, 20, 21,
                                        29, 12, 28, 17,
                                         1, 15, 23, 26,
                                         5, 18, 31, 10,
                                         2,  8, 24, 14,
                                        32, 27,  3,  9,
                                        19, 13, 30,  6,
                                        22, 11,  4, 25 );
    
    Constant Left_PC : PChoice_Table := ( 57, 49, 41, 33, 25, 17,  9,
                                           1, 58, 50, 42, 34, 26, 18,
                                          10,  2, 59, 51, 43, 35, 27,
                                          19, 11,  3, 60, 52, 44, 36 );

    Constant Right_PC : PChoice_Table := ( 63, 55, 47, 39, 31, 23, 15,
                                            7, 62, 54, 46, 38, 30, 22,
                                           14,  6, 61, 53, 45, 37, 29,
                                           21, 13,  5, 28, 20, 12,  4 );
    
    Constant Key_Permu : Permu_Sec_Table := ( 14, 17, 11, 24,  1,  5,
                                               3, 28, 15,  6, 21, 10,
                                              23, 19, 12,  4, 26,  8,
                                              16,  7, 27, 20, 13,  2,
                                              41, 52, 31, 37, 47, 55,
                                              30, 40, 51, 45, 33, 48,
                                              44, 49, 39, 56, 34, 53,
                                              46, 42, 50, 36, 29, 32 );
    
    Constant Sub_Box : S_Box := (
        ((14,4,13,1,2,15,11,8,3,10,6,12,5,9,0,7), -- S1
         (0,15,7,4,14,2,13,1,10,6,12,11,9,5,3,8),
         (4,1,14,8,13,6,2,11,15,12,9,7,3,10,5,0),
         (15,12,8,2,4,9,1,7,5,11,3,14,10,0,6,13)),
        ((15,1,8,14,6,11,3,4,9,7,2,13,12,0,5,10), -- S2
         (3,13,4,7,15,2,8,14,12,0,1,10,6,9,11,5),
         (0,14,7,11,10,4,13,1,5,8,12,6,9,3,2,15),
         (13,8,10,1,3,15,4,2,11,6,7,12,0,5,14,9)),
        ((10,0,9,14,6,3,15,5,1,13,12,7,11,4,2,8), -- S3
         (13,7,0,9,3,4,6,10,2,8,5,14,12,11,15,1),
         (13,6,4,9,8,15,3,0,11,1,2,12,5,10,14,7),
         (1,10,13,0,6,9,8,7,4,15,14,3,11,5,2,12)),
        ((7,13,14,3,0,6,9,10,1,2,8,5,11,12,4,15), -- S4
         (13,8,11,5,6,15,0,3,4,7,2,12,1,10,14,9),
         (10,6,9,0,12,11,7,13,15,1,3,14,5,2,8,4),
         (3,15,0,6,10,1,13,8,9,4,5,11,12,7,2,14)),
        ((2,12,4,1,7,10,11,6,8,5,3,15,13,0,14,9), -- S5
         (14,11,2,12,4,7,13,1,5,0,15,10,3,9,8,6),
         (4,2,1,11,10,13,7,8,15,9,12,5,6,3,0,14),
         (11,8,12,7,1,14,2,13,6,15,0,9,10,4,5,3)),
        ((12,1,10,15,9,2,6,8,0,13,3,4,14,7,5,11), -- S6
         (10,15,4,2,7,12,9,5,6,1,13,14,0,11,3,8),
         (9,14,15,5,2,8,12,3,7,0,4,10,1,13,11,6),
         (4,3,2,12,9,5,15,10,11,14,1,7,6,0,8,13)),
        ((4,11,2,14,15,0,8,13,3,12,9,7,5,10,6,1),  -- S7
         (13,0,11,7,4,9,1,10,14,3,5,12,2,15,8,6),
         (1,4,11,13,12,3,7,14,10,15,6,8,0,5,9,2),
         (6,11,13,8,1,4,10,7,9,5,0,15,14,2,3,12)),
        ((13,2,8,4,6,15,11,1,10,9,3,14,5,0,12,7), -- S8
         (1,15,13,8,10,3,7,4,12,5,6,11,0,14,9,2),
         (7,11,4,1,9,12,14,2,0,6,10,13,15,3,5,8),
         (2,1,14,7,4,10,8,13,15,12,9,0,3,5,6,11))
    );
    Constant Round_Shift : Shift_Table := ( 1, 1, 2, 2, 2, 2, 2, 2, 1, 2, 2, 2, 2, 2, 2, 1, 0 );

    -- Function Definition
    FUNCTION Permuation_Choice1( Signal Key : std_logic_vector; 
                                 Choice_Table : PChoice_Table ) RETURN std_logic_vector;
    
    FUNCTION Permuation_Choice2( Key : std_logic_vector;
                                 Choice_Table : Permu_Sec_Table ) RETURN std_logic_vector;
    
    FUNCTION Crypt_Process( Text : std_logic_vector;
                             Key : std_logic_vector ) RETURN std_logic_vector;
END PACKAGE DES_def;

PACKAGE BODY DES_def IS
    FUNCTION Permuation_Choice1( Signal Key : std_logic_vector;
                                 Choice_Table : PChoice_Table ) RETURN std_logic_vector IS
        Variable Choice_Key : std_logic_vector( 1 to 28 );
    BEGIN
        FOR I IN Choice_Key'left to Choice_Key'right LOOP
            Choice_Key(I) := Key(Choice_Table(I));
        END LOOP;
        RETURN Choice_Key;
    END Permuation_Choice1;

    FUNCTION Permuation_Choice2( Key : std_logic_vector;
                                 Choice_Table : Permu_Sec_Table) RETURN std_logic_vector IS
        Variable Choice_Key : std_logic_vector( 1 to 48 ) := (others => 'X');
    BEGIN
        FOR I IN Choice_Key'left to Choice_Key'right LOOP
            Choice_Key(I) := Key(Choice_Table(I));
        END LOOP;
        RETURN Choice_Key;
    END Permuation_Choice2;

    FUNCTION Crypt_Process( Text : std_logic_vector;  -- 32 downto 1
                             Key : std_logic_vector ) RETURN std_logic_vector IS
        Variable Temp_Text : std_logic_vector( 1 to 32 );
        Variable Result_Text : std_logic_vector( 1 to 32 );
        Variable Expan_Text : std_logic_vector( 1 to 48 );
        Variable row : std_logic_vector( 1 downto 0 );
        Variable col : std_logic_vector( 3 downto 0 );
    BEGIN
        -- Expand 32 bit to 48 bit
        FOR I IN 1 TO 48 LOOP
            Expan_Text(I) := Text( E_Table(I) );
        END LOOP;

        -- XOR with 48 bit key
        Expan_Text := Expan_Text XOR Key;

        -- Substitution Box
        FOR I IN 0 TO 7 LOOP
            row := Expan_Text( 1 + I * 6 ) & Expan_Text( 6 + I * 6 );
            col := Expan_Text( 2 + I * 6 ) & Expan_Text( 3 + I * 6 ) & Expan_Text( 4 + I * 6 ) & Expan_Text( 5 + I * 6 );
            Temp_Text( 1 + I * 4 to 4 + I * 4 ) := 
            std_logic_vector(to_unsigned(Sub_Box( I + 1 )( Conv_Integer(row), Conv_Integer(col)),4));
        END LOOP;

        -- Permutation
        FOR I IN 1 TO 32 LOOP
            Result_Text(I) := Temp_Text(P_Table(I));
        END LOOP;

        RETURN Result_Text;
    END Crypt_Process;
END PACKAGE BODY DES_def;

